module CU(
    input wire [5:0] opcode,
    output reg RegDest,
    output reg Jump,
    output reg Branch,
    output reg MemToReg,
    output reg [5:0] ALUOp,
    output reg MemWrite,
    output reg ALUsrc,
    output reg RegWrite,
    output reg jalCtrl,
    output reg jrCtrl
);


endmodule