`define INFINITY_POSITIVE_CONST 32'b01111111110000000000000000000000
`define INFINITY_NEGATIVE_CONST 32'b11111111110000000000000000000000
// https://stackoverflow.com/a/55648118
// https://en.wikipedia.org/wiki/NaN
`define QNAN_CONST 32'b?111111111??????????????????????
`define SNAN_CONST 32'b?111111110??????????????????????
