`define R_TYPE 6'b000000
`define J_TYPE 6'b00001?

// R Type macros


// J Type macros
`define J       6'b000010
`define JAL     6'b000011


// I Type macros
`define ADDi    6'b001000
`define ADDiu   6'b001001
`define ANDi    6'b001100
`define XORi    6'b001110
`define ORi     6'b001101
`define BEQ     6'b000100
`define BNE     6'b000101 
`define BLEZ    6'b000110 
`define BGTZ    6'b000111 
`define LW      6'b100011
`define SW      6'b101011
`define LB      6'b100000
`define SB      6'b101000
`define SLTi    6'b001010 





