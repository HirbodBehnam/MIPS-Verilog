`define R_TYPE 6'b000000
`define J_TYPE 6'b0000??

