`define FPU_ADD 4'b0000
`define FPU_SUB 4'b0001
`define FPU_MULT 4'b0010
`define FPU_DIV 4'b0011
`define FPU_NEGATE 4'b0100
`define FPU_ROUND 4'b0101
`define FPU_FLOAT_TO_BINARY 4'b0110
`define FPU_BINARY_TO_FLOAT 4'b0111
`define FPU_COMP_LT 4'b1000
`define FPU_COMP_LE 4'b1001
`define FPU_COMP_EQ 4'b1010
`define FPU_COMP_NQ 4'b1011
`define FPU_COMP_GT 4'b1100
`define FPU_COMP_GE 4'b1101
`define FPU_MOVE_TO_FLOAT 4'b1110
`define FPU_MOVE_TO_FLOAT 4'b1111