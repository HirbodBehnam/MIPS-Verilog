`define ALU_ADD 5'b00000
`define ALU_SUB 5'b00001
`define ALU_MULT 5'b00010
`define ALU_DIV 5'b00011

`define ALU_XOR 5'b00100
`define ALU_AND 5'b00101
`define ALU_OR 5'b00110
`define ALU_NOR 5'b00111

`define ALU_UNSIGNED_SHIFT_LEFT 5'b01000
`define ALU_UNSIGNED_SHIFT_RIGHT 5'b01001
`define ALU_UNSIGNED_SHIFT_LEFT_SH_AMOUNT 5'b01010
`define ALU_UNSIGNED_SHIFT_RIGHT_SH_AMOUNT 5'b01011
`define ALU_SIGNED_SHIFT_LEFT_SH_AMOUNT 5'b01100
`define ALU_SIGNED_SHIFT_RIGHT_SH_AMOUNT 5'b01101

`define ALU_COMP_GT 5'b10000
`define ALU_COMP_LT 5'b10001
`define ALU_COMP_GE 5'b10010
`define ALU_COMP_LE 5'b10011
`define ALU_COMP_EQ 5'b10100
`define ALU_COMP_NEQ 5'b10101

`define ALU_LUI 5'b11000