`include "fp_consts.sv";

module FP_Divider (
    input [31:0] a,
    input [31:0] b,
    output reg [31:0] result,
    output reg overflow,
    output reg underflow
);
    
endmodule