`define R_TYPE 6'b000000
`define J_TYPE 6'b00001?

// R Type macros


// J Type macros


// I Type macros
