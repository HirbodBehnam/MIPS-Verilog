module adder(output [31:0] res, input [31:0] a, input [31:0] b);
	assign res = a + b;
endmodule
