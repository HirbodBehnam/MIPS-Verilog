`define ALU_ADD 4'b0000
`define ALU_SUB 4'b0001
`define ALU_MULT 4'b0010
`define ALU_DIV 4'b0011

`define ALU_XOR 4'b0100
`define ALU_AND 4'b0101
`define ALU_OR 4'b0110
`define ALU_NOR 4'b0111

`define ALU_UNSIGNED_SHIFT_LEFT 4'b1000
`define ALU_UNSIGNED_SHIFT_RIGHT 4'b1001
`define ALU_SIGNED_SHIFT_LEFT 4'b1010
`define ALU_SIGNED_SHIFT_RIGHT 4'b1011

`define ALU_COMP_GT 4'b1100
`define ALU_COMP_LT 4'b1101
`define ALU_COMP_GE 4'b1110
`define ALU_ADD_LE 4'b1111