`define INFINITY_POSITIVE_CONST 32'b01111111100000000000000000000000
`define INFINITY_NEGATIVE_CONST 32'b11111111100000000000000000000000
// https://stackoverflow.com/a/55648118
// https://en.wikipedia.org/wiki/NaN
`define QNAN_CONST 32'b?111111111??????????????????????
`define SNAN_CONST 32'b?1111111101?????????????????????
`define QNAN_SAMPLE_CONST 32'b01111111110000000000000000000000
`define SNAN_SAMPLE_CONST 32'b01111111101000000000000000000000
`define ZERO 32'b00000000000000000000000000000000
// 0.5
`define POSITIVE_HALF 32'b00111111000000000000000000000000